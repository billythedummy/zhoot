package enemy_def;
    typedef enum {
        DEAD,
        ALIVE,
        DYING
    } enemy_state_t;
endpackage : enemy_def