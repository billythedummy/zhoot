module gunshot_player ();

endmodule