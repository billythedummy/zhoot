import enemy_def::*;

