module gunshot_rom (
    input logic clk,
    input logic [] addr,
    output logic [23:0] q
);
    

endmodule